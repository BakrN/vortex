
module VX_tensor_core#() () ;


endmodule;
