package tc_pkg;

    typedef enum logic[1:0] {
        ACC_SRC_ZERO = 2'b00,
        ACC_SRC_TILE,
        ACC_SRC_REG
    } acc_src_t;

endpackage
