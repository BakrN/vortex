module pe_group #() (


    );

    // Signals shared across all PEs
    logic wid;
    logic wb ;
    logic rd ; // These will be shared have to
    // can change after FPU Latency


endmodule
